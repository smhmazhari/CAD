module ();
checker_top_module  #(
    parameter IF_CELL_SIZE = 8 ,
    parameter IF_ADDRESS_SIZE = 8 ,
    parameter FILTER_CELL_SIZE = 8 ,
    parameter FILTER_ADDRESS_SIZE = 8 ,
    parameter STRIDE_SIZE = 2 ,
    parameter CELL_NUMS_IF = 8,
    parameter CELL_NUMS_FILTER = 8  
)(
          input clk,
          input rst,
          input inner_start,
          input [STRIDE_SIZE:0] stride,
          input [2:0] filter_size,
          input [2:0] if_size,
          input write_cnt_if,
          input write_cnt_filter,
          input [IF_ADDRESS_SIZE:0] write_addr_if,
          input [FILTER_ADDRESS_SIZE:0] write_addr_filter,
          output scratch_write_en,
          output par_done,
          output can_count,
          output can_mult,
          output Done
    
);

endmodule