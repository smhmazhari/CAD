module shift_register_left_16bit (
  input clk,  
  input load,
  input shl, 
  input [15:0] data_in, 
  output[15:0] data_out 
);


  shift_block b15(clk,rst,load,shl,data_in[15],data_out[14],data_out[15]);
  shift_block b14(clk,rst,load,shl,data_in[14],data_out[13],data_out[14]);
  shift_block b13(clk,rst,load,shl,data_in[13],data_out[12],data_out[13]);
  shift_block b12(clk,rst,load,shl,data_in[12],data_out[11],data_out[12]);
  shift_block b11(clk,rst,load,shl,data_in[11],data_out[10],data_out[11]);
  shift_block b10(clk,rst,load,shl,data_in[10],data_out[9],data_out[10]);
  shift_block b9(clk,rst,load,shl,data_in[9],data_out[8],data_out[9]);
  shift_block b8(clk,rst,load,shl,data_in[8],data_out[7],data_out[8]);
  shift_block b7(clk,rst,load,shl,data_in[7],data_out[6],data_out[7]);
  shift_block b6(clk,rst,load,shl,data_in[6],data_out[5],data_out[6]);
  shift_block b5(clk,rst,load,shl,data_in[5],data_out[4],data_out[5]);
  shift_block b4(clk,rst,load,shl,data_in[4],data_out[3],data_out[4]);
  shift_block b3(clk,rst,load,shl,data_in[3],data_out[2],data_out[3]);
  shift_block b2(clk,rst,load,shl,data_in[2],data_out[1],data_out[2]);
  shift_block b1(clk,rst,load,shl,data_in[1],data_out[0],data_out[1]);
  shift_block b0(clk,rst,load,shl,data_in[0],1'd0,data_out[0]);
endmodule